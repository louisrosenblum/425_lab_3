*****************************************************************************
* CDL Netlist:
* Cell Name: and2
* Netlisted on: Apr 21 15:50:52 2022
*****************************************************************************


*****************************************************************************
* Global Net Declarations
*****************************************************************************
*.GLOBAL vdd! gnd!


*****************************************************************************
* PIN Control Statement
*****************************************************************************
*.PIN vdd! gnd!


*****************************************************************************
* BIPOLAR Declarations
*****************************************************************************
*.BIPOLAR
*.RESI = 2000.000000
*.SCALE METER


*****************************************************************************
* Parameter Statement
*****************************************************************************
.PARAM


*******************************************************************************
* Main Circuit Netlist:                                                       *
*                                                                             *
* Library: Lab4                                                               *
* Cell   : and2                                                               *
* View   : schematic                                                          *
* Last Time Saved: Apr 21 15:43:33 2022                                       *
*******************************************************************************
.subckt and2 F A B
*.PININFO F:O A:I B:I 
.ends and2
