*****************************************************************************
* CDL Netlist:
* Cell Name: four_bit_adder
* Netlisted on: Apr 23 00:22:59 2022
*****************************************************************************


*****************************************************************************
* Global Net Declarations
*****************************************************************************
*.GLOBAL vdd! gnd!


*****************************************************************************
* PIN Control Statement
*****************************************************************************
*.PIN vdd! gnd!


*****************************************************************************
* BIPOLAR Declarations
*****************************************************************************
*.BIPOLAR
*.RESI = 2000.000000
*.SCALE METER


*****************************************************************************
* Parameter Statement
*****************************************************************************
.PARAM


*******************************************************************************
* Sub-Circuit Netlist:                                                        *
*                                                                             *
* Library: Lab4                                                               *
* Cell   : one_bit_adder                                                      *
* View   : schematic                                                          *
* Last Time Saved: Apr  3 20:56:03 2022                                       *
*******************************************************************************
.subckt one_bit_adder Cout Sum A B Cin
*.PININFO Cout:O Sum:O A:I B:I Cin:I 
.ends one_bit_adder


*******************************************************************************
* Main Circuit Netlist:                                                       *
*                                                                             *
* Library: Lab4                                                               *
* Cell   : four_bit_adder                                                     *
* View   : schematic                                                          *
* Last Time Saved: Apr 22 22:31:20 2022                                       *
*******************************************************************************
.subckt four_bit_adder Cout Sum0 Sum1 Sum2 Sum3 A0 A1 A2 A3 B0 B1 B2 B3
*.PININFO Cout:O Sum0:O Sum1:O Sum2:O Sum3:O A0:I A1:I A2:I A3:I B0:I B1:I B2:I
*.PININFO B3:I 
XI3 Cout Sum3 A3 B3 net35 one_bit_adder
XI2 net35 Sum2 A2 B2 net030 one_bit_adder
XI1 net030 Sum1 A1 B1 net033 one_bit_adder
XI0 net033 Sum0 A0 B0 gnd! one_bit_adder
.ends four_bit_adder
