*****************************************************************************
* CDL Netlist:
* Cell Name: or3
* Netlisted on: Apr 25 10:33:43 2022
*****************************************************************************


*****************************************************************************
* Global Net Declarations
*****************************************************************************
*.GLOBAL vdd! gnd!


*****************************************************************************
* PIN Control Statement
*****************************************************************************
*.PIN vdd! gnd!


*****************************************************************************
* BIPOLAR Declarations
*****************************************************************************
*.BIPOLAR
*.RESI = 2000.000000
*.SCALE METER


*****************************************************************************
* Parameter Statement
*****************************************************************************
.PARAM


*******************************************************************************
* Sub-Circuit Netlist:                                                        *
*                                                                             *
* Library: Lab4                                                               *
* Cell   : or3                                                                *
* View   : schematic                                                          *
* Last Time Saved: Apr 22 21:36:12 2022                                       *
*******************************************************************************
.subckt or3 F A B C
*.PININFO F:O A:I B:I C:I 
.ends or3
