*****************************************************************************
* CDL Netlist:
* Cell Name: one_bit_adder_Leg3
* Netlisted on: Apr  3 20:24:21 2022
*****************************************************************************


*****************************************************************************
* Global Net Declarations
*****************************************************************************
*.GLOBAL vdd! gnd!


*****************************************************************************
* PIN Control Statement
*****************************************************************************
*.PIN vdd! gnd!


*****************************************************************************
* BIPOLAR Declarations
*****************************************************************************
*.BIPOLAR
*.RESI = 2000.000000
*.SCALE METER


*****************************************************************************
* Parameter Statement
*****************************************************************************
.PARAM


*******************************************************************************
* Main Circuit Netlist:                                                       *
*                                                                             *
* Library: Lab4                                                               *
* Cell   : one_bit_adder_Leg3                                                 *
* View   : schematic                                                          *
* Last Time Saved: Apr  3 20:13:54 2022                                       *
*******************************************************************************
.subckt one_bit_adder_Leg3 Cout SumNot A B Cin
*.PININFO Cout:O SumNot:O A:I B:I Cin:I 
.ends one_bit_adder_Leg3
