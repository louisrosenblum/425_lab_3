*****************************************************************************
* CDL Netlist:
* Cell Name: d_flip_flop
* Netlisted on: Apr 23 00:46:42 2022
*****************************************************************************


*****************************************************************************
* Global Net Declarations
*****************************************************************************
*.GLOBAL vdd! gnd!


*****************************************************************************
* PIN Control Statement
*****************************************************************************
*.PIN vdd! gnd!


*****************************************************************************
* BIPOLAR Declarations
*****************************************************************************
*.BIPOLAR
*.RESI = 2000.000000
*.SCALE METER


*****************************************************************************
* Parameter Statement
*****************************************************************************
.PARAM


*******************************************************************************
* Sub-Circuit Netlist:                                                        *
*                                                                             *
* Library: Lab4                                                               *
* Cell   : d_flip_flop                                                        *
* View   : schematic                                                          *
* Last Time Saved: Apr 10 02:58:43 2022                                       *
*******************************************************************************
.subckt d_flip_flop Q Clk D
*.PININFO Q:O Clk:I D:I 
.ends d_flip_flop
