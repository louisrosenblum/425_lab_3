*****************************************************************************
* CDL Netlist:
* Cell Name: one_bit_adder_Leg1
* Netlisted on: Apr  3 14:27:40 2022
*****************************************************************************


*****************************************************************************
* Global Net Declarations
*****************************************************************************
*.GLOBAL gnd! vdd!


*****************************************************************************
* PIN Control Statement
*****************************************************************************
*.PIN gnd! vdd!


*****************************************************************************
* BIPOLAR Declarations
*****************************************************************************
*.BIPOLAR
*.RESI = 2000.000000
*.SCALE METER


*****************************************************************************
* Parameter Statement
*****************************************************************************
.PARAM


*******************************************************************************
* Main Circuit Netlist:                                                       *
*                                                                             *
* Library: Lab4                                                               *
* Cell   : one_bit_adder_Leg1                                                 *
* View   : schematic                                                          *
* Last Time Saved: Apr  3 11:30:04 2022                                       *
*******************************************************************************
.subckt one_bit_adder_Leg1 CoutNot A B Cin
*.PININFO CoutNot:O A:I B:I Cin:I 
.ends one_bit_adder_Leg1
