*****************************************************************************
* CDL Netlist:
* Cell Name: one_bit_adder_Leg4
* Netlisted on: Apr  3 22:11:02 2022
*****************************************************************************


*****************************************************************************
* Global Net Declarations
*****************************************************************************
*.GLOBAL gnd! vdd!


*****************************************************************************
* PIN Control Statement
*****************************************************************************
*.PIN gnd! vdd!


*****************************************************************************
* BIPOLAR Declarations
*****************************************************************************
*.BIPOLAR
*.RESI = 2000.000000
*.SCALE METER


*****************************************************************************
* Parameter Statement
*****************************************************************************
.PARAM


*******************************************************************************
* Main Circuit Netlist:                                                       *
*                                                                             *
* Library: Lab4                                                               *
* Cell   : one_bit_adder_Leg4                                                 *
* View   : schematic                                                          *
* Last Time Saved: Apr  3 20:56:03 2022                                       *
*******************************************************************************
.subckt one_bit_adder_Leg4 Cout Sum A B Cin
*.PININFO Cout:O Sum:O A:I B:I Cin:I 
.ends one_bit_adder_Leg4
